module fetch_unit(input clk,rst
