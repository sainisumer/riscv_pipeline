module fetch_unit
